module decoder(input logic [4:0]sel, output logic [31:0]Y);

always_comb begin
		case(sel)
			5'd0:  Y = 32'b00000000000000000000000000000001;
			5'd1:  Y = 32'b00000000000000000000000000000010;
			5'd2:  Y = 32'b00000000000000000000000000000100;
			5'd3:  Y = 32'b00000000000000000000000000001000;
			5'd4:  Y = 32'b00000000000000000000000000010000;
			5'd5:  Y = 32'b00000000000000000000000000100000;
			5'd6:  Y = 32'b00000000000000000000000001000000;
			5'd7:  Y = 32'b00000000000000000000000010000000;
			5'd8:  Y = 32'b00000000000000000000000100000000;
			5'd9:  Y = 32'b00000000000000000000001000000000;
			5'd10: Y = 32'b00000000000000000000010000000000;
			5'd11: Y = 32'b00000000000000000000100000000000;
			5'd12: Y = 32'b00000000000000000001000000000000;
			5'd13: Y = 32'b00000000000000000010000000000000;
			5'd14: Y = 32'b00000000000000000100000000000000;
			5'd15: Y = 32'b00000000000000001000000000000000;
			5'd16: Y = 32'b00000000000000010000000000000000;
			5'd17: Y = 32'b00000000000000100000000000000000;
			5'd18: Y = 32'b00000000000001000000000000000000;
			5'd19: Y = 32'b00000000000010000000000000000000;
			5'd20: Y = 32'b00000000000100000000000000000000;
			5'd21: Y = 32'b00000000001000000000000000000000;
			5'd22: Y = 32'b00000000010000000000000000000000;
			5'd23: Y = 32'b00000000100000000000000000000000;
			5'd24: Y = 32'b00000001000000000000000000000000;
			5'd25: Y = 32'b00000010000000000000000000000000;
			5'd26: Y = 32'b00000100000000000000000000000000;
			5'd27: Y = 32'b00001000000000000000000000000000;
			5'd28: Y = 32'b00010000000000000000000000000000;
			5'd29: Y = 32'b00100000000000000000000000000000;
			5'd30: Y = 32'b01000000000000000000000000000000;
			5'd31: Y = 32'b10000000000000000000000000000000;
		endcase
	end
endmodule
