library verilog;
use verilog.vl_types.all;
entity flopenr_tb is
end flopenr_tb;
