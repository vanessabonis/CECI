library verilog;
use verilog.vl_types.all;
entity flopr_tb is
end flopr_tb;
