library verilog;
use verilog.vl_types.all;
entity bancoRegistradores_tb is
end bancoRegistradores_tb;
