library verilog;
use verilog.vl_types.all;
entity decoder_tb is
end decoder_tb;
