library verilog;
use verilog.vl_types.all;
entity mux2_tb is
end mux2_tb;
