library verilog;
use verilog.vl_types.all;
entity ShiftPC_tb is
end ShiftPC_tb;
