library verilog;
use verilog.vl_types.all;
entity SignExtend_tb is
end SignExtend_tb;
