library verilog;
use verilog.vl_types.all;
entity inversor is
    port(
        a               : in     vl_logic;
        y               : out    vl_logic
    );
end inversor;
