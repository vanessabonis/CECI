library verilog;
use verilog.vl_types.all;
entity mux4_tb is
end mux4_tb;
