library verilog;
use verilog.vl_types.all;
entity ShiftLeft2_tb is
end ShiftLeft2_tb;
