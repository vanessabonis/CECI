library verilog;
use verilog.vl_types.all;
entity ULA_1bit_tb is
end ULA_1bit_tb;
